module teste(input a, output b);
    assign b = a;
endmodule